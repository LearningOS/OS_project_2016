-------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
-------------------------------------------------------------------------------------
package defines is
-------------------------------------------------------------------------------------

	type regs32 is array (31 downto 0) of std_logic_vector(31 downto 0);
	type brk_arr is array (3 downto 0) of std_logic_vector(32 downto 0);
	type wtc_arr is array (3 downto 0) of std_logic_vector(33 downto 0);
	--type type_digit7 is array (6 downto 0) of std_logic_vector;

	
-------------------------------------------------------------------------------------
end package;

package body defines is
-------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------
end defines;
-------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------